module u_lsu (
input clk,
input rstn,
// input
input        lsu_e,
input        lsu_w,
input [31:0] lsu_a,

);


